** sch_path: /foss/designs/tt10-uR-IPs/xschem/MND_ES-4.sch
**.subckt MND_ES-4
XM2 vds vgs GND GND sky130_fd_pr__nfet_01v8 L=2 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
vs_vgs vgs GND 1.8
.save i(vs_vgs)
vs_vds vds GND 1.8
.save i(vs_vds)
**** begin user architecture code


.option gmin=1e-12


.dc vs_vgs 0 5 0.01 vs_vds 0 5 0.5

.save all
*write es4.raw




** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
