magic
tech sky130A
magscale 1 2
timestamp 1741544095
<< locali >>
rect 27845 1407 27879 1722
<< viali >>
rect 27845 1373 27879 1407
<< metal1 >>
rect 27715 2498 27743 2864
rect 26598 2470 27743 2498
rect 26598 2309 26626 2470
rect 29942 2251 30525 2299
rect 26235 2126 26299 2132
rect 26235 2074 26241 2126
rect 26293 2114 26299 2126
rect 26293 2086 26555 2114
rect 26293 2074 26299 2086
rect 26235 2068 26299 2074
rect 27126 1968 27178 1974
rect 27126 1910 27178 1916
rect 27725 1663 27777 1669
rect 27725 1605 27777 1611
rect 28326 1663 28378 1669
rect 28326 1605 28378 1611
rect 28881 1663 28933 1669
rect 28881 1605 28933 1611
rect 29436 1663 29488 1669
rect 29436 1605 29488 1611
rect 28893 1604 28921 1605
rect 30477 1462 30525 2251
rect 30477 1416 30526 1462
rect 27833 1407 27891 1413
rect 27833 1373 27845 1407
rect 27879 1373 27891 1407
rect 27833 1367 27891 1373
rect 26498 1077 26678 1078
rect 27845 1077 27879 1367
rect 30478 1356 30526 1416
rect 26498 1043 27879 1077
rect 30477 1336 30526 1356
rect 26498 894 26678 1043
rect 30477 984 30525 1336
rect 26492 714 26498 894
rect 26678 714 26684 894
rect 30362 732 30542 984
rect 30356 552 30362 732
rect 30542 552 30548 732
<< via1 >>
rect 26241 2074 26293 2126
rect 27126 1916 27178 1968
rect 27725 1611 27777 1663
rect 28326 1611 28378 1663
rect 28881 1611 28933 1663
rect 29436 1611 29488 1663
rect 26498 714 26678 894
rect 30362 552 30542 732
<< metal2 >>
rect 26175 2617 27749 2645
rect 26175 2137 26203 2617
rect 27074 2157 27254 2185
rect 26161 2132 26235 2137
rect 26161 2128 26299 2132
rect 26161 2072 26170 2128
rect 26226 2126 26299 2128
rect 26226 2074 26241 2126
rect 26293 2074 26299 2126
rect 26226 2072 26299 2074
rect 26161 2068 26299 2072
rect 26161 2063 26235 2068
rect 27011 1912 27020 1968
rect 27076 1954 27085 1968
rect 27120 1954 27126 1968
rect 27076 1926 27126 1954
rect 27076 1912 27085 1926
rect 27120 1916 27126 1926
rect 27178 1916 27184 1968
rect 27226 1651 27254 2157
rect 27282 1912 27291 1968
rect 27347 1954 27356 1968
rect 27347 1926 27743 1954
rect 27347 1912 27356 1926
rect 27719 1651 27725 1663
rect 27226 1623 27725 1651
rect 27719 1611 27725 1623
rect 27777 1611 27783 1663
rect 28320 1611 28326 1663
rect 28378 1611 28384 1663
rect 28875 1611 28881 1663
rect 28933 1611 28939 1663
rect 29430 1611 29436 1663
rect 29488 1654 29494 1663
rect 29488 1620 29720 1654
rect 29488 1611 29494 1620
rect 28338 1428 28366 1611
rect 28875 1605 28939 1611
rect 28893 1428 28921 1605
rect 29692 1428 29720 1620
rect 28315 1372 28324 1428
rect 28380 1372 28389 1428
rect 28870 1372 28879 1428
rect 28935 1372 28944 1428
rect 29669 1372 29678 1428
rect 29734 1372 29743 1428
rect 26498 894 26678 900
rect 26498 527 26678 714
rect 30362 732 30542 738
rect 26494 357 26503 527
rect 26673 357 26682 527
rect 30362 519 30542 552
rect 26498 352 26678 357
rect 30358 349 30367 519
rect 30537 349 30546 519
rect 30362 344 30542 349
<< via2 >>
rect 26170 2072 26226 2128
rect 27020 1912 27076 1968
rect 27291 1912 27347 1968
rect 28324 1372 28380 1428
rect 28879 1372 28935 1428
rect 29678 1372 29734 1428
rect 26503 357 26673 527
rect 30367 349 30537 519
<< metal3 >>
rect 370 2131 446 2137
rect 370 2067 376 2131
rect 440 2130 446 2131
rect 26161 2130 26231 2133
rect 440 2128 26231 2130
rect 440 2072 26170 2128
rect 26226 2072 26231 2128
rect 440 2070 26231 2072
rect 440 2067 446 2070
rect 26161 2067 26231 2070
rect 370 2061 446 2067
rect 26092 1908 26098 1972
rect 26162 1970 26168 1972
rect 27015 1970 27081 1973
rect 27286 1970 27352 1973
rect 26162 1968 27352 1970
rect 26162 1912 27020 1968
rect 27076 1912 27291 1968
rect 27347 1912 27352 1968
rect 26162 1910 27352 1912
rect 26162 1908 26168 1910
rect 27015 1907 27081 1910
rect 27286 1907 27352 1910
rect 28322 1433 28382 1742
rect 28877 1433 28937 1733
rect 29676 1433 29736 1757
rect 28319 1428 28385 1433
rect 28319 1372 28324 1428
rect 28380 1372 28385 1428
rect 28319 1367 28385 1372
rect 28874 1428 28940 1433
rect 28874 1372 28879 1428
rect 28935 1372 28940 1428
rect 28874 1367 28940 1372
rect 29673 1428 29739 1433
rect 29673 1372 29678 1428
rect 29734 1372 29739 1428
rect 29673 1367 29739 1372
rect 26498 527 26678 532
rect 26498 357 26503 527
rect 26673 357 26678 527
rect 26498 199 26678 357
rect 30362 519 30542 524
rect 30362 349 30367 519
rect 30537 349 30542 519
rect 30362 199 30542 349
rect 26493 21 26499 199
rect 26677 21 26683 199
rect 30357 21 30363 199
rect 30541 21 30547 199
rect 26498 20 26678 21
rect 30362 20 30542 21
<< via3 >>
rect 376 2067 440 2131
rect 26098 1908 26162 1972
rect 26499 21 26677 199
rect 30363 21 30541 199
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 2131 600 44152
rect 200 2067 376 2131
rect 440 2067 600 2131
rect 200 1000 600 2067
rect 800 1970 1200 44152
rect 26097 2663 30085 2723
rect 26097 2662 27784 2663
rect 26097 1973 26158 2662
rect 26097 1972 26163 1973
rect 26097 1970 26098 1972
rect 800 1910 26098 1970
rect 800 1000 1200 1910
rect 26097 1908 26098 1910
rect 26162 1908 26163 1972
rect 26097 1907 26163 1908
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 199 26678 200
rect 26498 21 26499 199
rect 26677 21 26678 199
rect 26498 0 26678 21
rect 30362 199 30542 200
rect 30362 21 30363 199
rect 30541 21 30542 199
rect 30362 0 30542 21
use ibias_10nA  bias /foss/designs/tt10-uR-IPs/magic/tt10/biasGen
timestamp 1741542799
transform 1 0 26376 0 1 3242
box 108 -1612 850 -889
use osc  osc_0 /foss/designs/tt10-uR-IPs/magic/tt10/osc
timestamp 1741541561
transform 1 0 27735 0 1 1603
box -20 1 2272 1261
use s130_mim_dl_40fF  cap_osc_1 /foss/designs/tt10-uR-IPs/magic/tt10/osc/cap
timestamp 1741537464
transform -1 0 29612 0 -1 2002
box -597 -828 59 329
use s130_mim_dl_40fF  cap_osc_2 /foss/designs/tt10-uR-IPs/magic/tt10/osc/cap
timestamp 1741537464
transform -1 0 27820 0 -1 2002
box -597 -828 59 329
use s130_mim_dl_40fF  cap_osc_3 /foss/designs/tt10-uR-IPs/magic/tt10/osc/cap
timestamp 1741537464
transform -1 0 28716 0 -1 2002
box -597 -828 59 329
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
