** sch_path: /foss/designs/tt10-uR-IPs/xschem/schmitt_trigger_ro.sch
.subckt schmitt_trigger_ro Vdd Vin Vout Vss
*.PININFO Vdd:I Vss:I Vin:I Vout:O
XM10 net1 Vin Vdd Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=1 m=1
XM2 Vout Vin net1 Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=1 m=1
XM4 net3 Vout net1 Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=1 m=1
XM6 Vout Vin net2 Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
XM1 net2 Vin Vss Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
XM3 Vdd Vout net2 Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
.ends
.end
