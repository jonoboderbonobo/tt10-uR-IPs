magic
tech sky130A
timestamp 1738500547
<< checkpaint >>
rect -649 -654 971 926
use sky130_fd_sc_hd__xnor2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 0 0 1 0
box -19 -24 341 296
<< end >>
