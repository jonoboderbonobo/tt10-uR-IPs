** sch_path: /foss/designs/tt10-uR-IPs/xschem/relax_osc_tb.sch
**.subckt relax_osc_tb
V2 vdd_hi GND 1.8
C1 net1 GND 10f m=1
.save v(vdd_hi)
.save v(out)
x1 vdd_hi out GND relax_osc
**** begin user architecture code


.control
*set filetype=ascii
*save all

op
tran 0.1n 1u

write tb_inv.raw
*exit

.endc



** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  relax_osc.sym # of pins=3
** sym_path: /foss/designs/tt10-uR-IPs/xschem/relax_osc.sym
** sch_path: /foss/designs/tt10-uR-IPs/xschem/relax_osc.sch
.subckt relax_osc Vdd Vout Vss
*.ipin Vss
*.ipin Vdd
*.opin Vout
R1 net1 Vout sky130_fd_pr__res_generic_l1 W=1 L=3000 m=1
XC1 net1 Vss sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=1 m=1
x1 Vdd net1 Vout Vss schmitt_trigger_ro
.ends


* expanding   symbol:  schmitt_trigger_ro.sym # of pins=4
** sym_path: /foss/designs/tt10-uR-IPs/xschem/schmitt_trigger_ro.sym
** sch_path: /foss/designs/tt10-uR-IPs/xschem/schmitt_trigger_ro.sch
.subckt schmitt_trigger_ro Vdd Vin Vout Vss
*.ipin Vdd
*.ipin Vss
*.ipin Vin
*.opin Vout
XM10 net1 Vin Vdd Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin net1 Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 Vout net1 Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout Vin net2 Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 Vin Vss Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vdd Vout net2 Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
