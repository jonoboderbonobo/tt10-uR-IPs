** sch_path: /foss/designs/tt10-uR-IPs/xschem/relax_osc.sch
**.subckt relax_osc Vdd Vout Vss
*.ipin Vss
*.ipin Vdd
*.opin Vout
R1 net1 Vout sky130_fd_pr__res_generic_l1 W=1 L=3000 m=1
XC1 net1 Vss sky130_fd_pr__cap_mim_m3_1 W=100 L=100 MF=1 m=1
x1 Vdd net1 Vout Vss schmitt_trigger_ro
**.ends
.end
