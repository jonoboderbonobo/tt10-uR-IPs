magic
tech sky130A
magscale 1 2
timestamp 1741560675
<< nwell >>
rect 934 -842 1557 -818
rect 934 -847 1234 -842
rect 1143 -851 1234 -847
rect 1152 -894 1234 -851
rect 1315 -847 1557 -842
rect 1315 -894 1453 -847
rect 1478 -894 1557 -847
rect 1152 -895 1291 -894
rect 1315 -895 1557 -894
rect 1152 -997 1557 -895
rect 1064 -1056 1104 -1050
rect 1064 -1077 1110 -1056
rect 1145 -1072 1557 -997
rect 1145 -1074 1239 -1072
rect 1145 -1082 1223 -1074
rect 1284 -1184 1557 -1072
rect 1230 -1365 1557 -1184
rect 1315 -1387 1483 -1365
<< psubdiff >>
rect 1297 -2106 1443 -2094
rect 1286 -2140 1310 -2106
rect 1432 -2140 1456 -2106
rect 1297 -2152 1443 -2140
<< nsubdiff >>
rect 1339 -1205 1446 -1193
rect 1328 -1239 1352 -1205
rect 1432 -1239 1456 -1205
rect 1339 -1251 1446 -1239
<< psubdiffcont >>
rect 1310 -2140 1432 -2106
<< nsubdiffcont >>
rect 1352 -1239 1432 -1205
<< poly >>
rect 1028 -1129 1058 -1075
rect 1028 -1376 1058 -1329
rect 1115 -1359 1145 -1329
rect 934 -1410 1058 -1376
rect 1028 -1422 1058 -1410
rect 1100 -1376 1165 -1359
rect 1378 -1376 1443 -1360
rect 1100 -1410 1115 -1376
rect 1149 -1410 1393 -1376
rect 1427 -1410 1443 -1376
rect 1100 -1426 1165 -1410
rect 1378 -1426 1443 -1410
rect 1115 -1448 1145 -1426
rect 1028 -1703 1058 -1648
<< polycont >>
rect 1115 -1410 1149 -1376
rect 1393 -1410 1427 -1376
<< locali >>
rect 982 -837 1172 -803
rect 982 -904 1016 -837
rect 1138 -931 1172 -837
rect 1138 -965 1303 -931
rect 1328 -1239 1352 -1205
rect 1432 -1239 1456 -1205
rect 982 -1333 1010 -1299
rect 1157 -1333 1303 -1299
rect 982 -1376 1016 -1333
rect 982 -1410 1115 -1376
rect 1149 -1410 1165 -1376
rect 982 -1444 1016 -1410
rect 982 -1478 1010 -1444
rect 1269 -1521 1303 -1333
rect 1377 -1410 1393 -1376
rect 1427 -1410 1443 -1376
rect 982 -1945 1016 -1903
rect 982 -1979 1270 -1945
rect 1286 -2140 1310 -2106
rect 1432 -2140 1456 -2106
<< viali >>
rect 1352 -1239 1432 -1205
rect 1115 -1410 1149 -1376
rect 1393 -1410 1427 -1376
rect 1310 -2140 1432 -2106
<< metal1 >>
rect 1315 -894 1381 -839
rect 1409 -950 1437 -935
rect 1064 -1056 1104 -1050
rect 1064 -1129 1110 -1056
rect 1269 -1193 1303 -1129
rect 1100 -1370 1165 -1369
rect 1100 -1376 1171 -1370
rect 1100 -1410 1115 -1376
rect 1149 -1410 1171 -1376
rect 1100 -1416 1171 -1410
rect 1268 -1448 1303 -1193
rect 1400 -1199 1428 -1087
rect 1346 -1205 1444 -1199
rect 1340 -1239 1352 -1205
rect 1432 -1239 1444 -1205
rect 1346 -1245 1444 -1239
rect 1378 -1376 1449 -1369
rect 1378 -1410 1393 -1376
rect 1427 -1410 1449 -1376
rect 1378 -1416 1449 -1410
rect 1151 -1486 1303 -1448
rect 1151 -1494 1197 -1486
rect 1064 -1702 1110 -1648
rect 1419 -1933 1447 -1929
rect 1410 -1975 1447 -1933
rect 1277 -2053 1349 -2007
rect 1410 -2100 1438 -1975
rect 1304 -2106 1438 -2100
rect 1298 -2140 1310 -2106
rect 1432 -2140 1444 -2106
rect 1304 -2146 1438 -2140
use sky130_fd_pr__nfet_01v8_QRJQW7  M1
timestamp 1741556153
transform 1 0 1130 0 1 -1548
box -65 -126 73 126
use sky130_fd_pr__nfet_01v8_2SPF2Z  M2
timestamp 1741556153
transform 1 0 1043 0 1 -1802
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_2JZFD3  M3
timestamp 1741556153
transform 1 0 1043 0 1 -1517
box -73 -157 73 95
use sky130_fd_pr__pfet_01v8_EJJ636_2  M4
timestamp 1741556153
transform 1 0 1130 0 1 -1229
box -65 -136 153 162
use sky130_fd_pr__pfet_01v8_EJJ636  M5
timestamp 1741556153
transform 1 0 1043 0 1 -1229
box -109 -136 109 162
use sky130_fd_pr__pfet_01v8_WXG636  M6
timestamp 1741556153
transform 1 0 1043 0 1 -975
box -109 -136 109 136
use sky130_fd_pr__nfet_01v8_3RATTY  M88
timestamp 1741560270
transform 1 0 1355 0 1 -1781
box -98 -282 98 282
use sky130_fd_pr__pfet_01v8_HW9MHL  M99
timestamp 1741556153
transform 1 0 1350 0 1 -999
box -129 -198 129 160
<< end >>
