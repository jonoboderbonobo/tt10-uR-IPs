magic
tech sky130A
magscale 1 2
timestamp 1738528573
<< viali >>
rect 6288 43847 6322 43881
rect 6515 43847 6549 43881
rect 6661 43726 6695 43760
<< metal1 >>
rect 6086 44223 6117 44224
rect 5815 44221 6117 44223
rect 1984 44196 6117 44221
rect 1984 44194 6088 44196
rect 1984 44193 6030 44194
rect 1787 44091 1793 44143
rect 1845 44133 1851 44143
rect 1984 44133 2012 44193
rect 5815 44192 6030 44193
rect 1845 44100 2015 44133
rect 1845 44091 1851 44100
rect 5795 43896 5857 43902
rect 7027 43900 7097 43906
rect 5795 43891 6338 43896
rect 5795 43839 5800 43891
rect 5852 43881 6338 43891
rect 5852 43847 6288 43881
rect 6322 43847 6338 43881
rect 5852 43839 6338 43847
rect 5795 43836 6338 43839
rect 6500 43891 7097 43900
rect 6500 43881 7036 43891
rect 6500 43847 6515 43881
rect 6549 43847 7036 43881
rect 6500 43839 7036 43847
rect 7088 43839 7097 43891
rect 5795 43834 6300 43836
rect 5795 43828 5857 43834
rect 6500 43830 7097 43839
rect 7027 43824 7097 43830
rect 6642 43779 6800 43780
rect 7271 43779 7337 43785
rect 6642 43772 7337 43779
rect 6642 43760 7278 43772
rect 6642 43726 6661 43760
rect 6695 43726 7278 43760
rect 6642 43720 7278 43726
rect 7330 43720 7337 43772
rect 6642 43713 7337 43720
rect 6642 43712 6800 43713
rect 7271 43707 7337 43713
rect 4463 43574 4469 43626
rect 4521 43615 4527 43626
rect 4521 43584 6126 43615
rect 4521 43574 4527 43584
<< via1 >>
rect 1793 44091 1845 44143
rect 5800 43839 5852 43891
rect 7036 43839 7088 43891
rect 7278 43720 7330 43772
rect 4469 43574 4521 43626
<< metal2 >>
rect 19941 44779 20003 44788
rect 5795 44723 19941 44779
rect 20003 44723 20053 44779
rect 5795 44717 20053 44723
rect 1632 44090 1641 44146
rect 1697 44134 1706 44146
rect 1793 44143 1845 44149
rect 1697 44101 1793 44134
rect 1697 44090 1706 44101
rect 1793 44085 1845 44091
rect 5795 43896 5857 44717
rect 19941 44714 20003 44717
rect 7027 44637 7097 44638
rect 7027 44567 19365 44637
rect 19435 44567 19457 44637
rect 7027 43900 7097 44567
rect 18843 44342 18909 44351
rect 7271 44286 18843 44342
rect 7271 44276 18909 44286
rect 5789 43891 5863 43896
rect 5789 43839 5800 43891
rect 5852 43839 5863 43891
rect 5789 43834 5863 43839
rect 7021 43891 7103 43900
rect 7021 43839 7036 43891
rect 7088 43839 7103 43891
rect 7021 43830 7103 43839
rect 7271 43779 7337 44276
rect 7265 43772 7343 43779
rect 7265 43720 7278 43772
rect 7330 43720 7343 43772
rect 7265 43713 7343 43720
rect 4263 43629 4319 43638
rect 4469 43626 4521 43632
rect 4319 43585 4469 43616
rect 4263 43564 4319 43573
rect 4469 43568 4521 43574
<< via2 >>
rect 19941 44723 20003 44779
rect 1641 44090 1697 44146
rect 19365 44567 19435 44637
rect 18843 44286 18909 44342
rect 4263 43573 4319 43629
<< metal3 >>
rect 18843 45027 18909 45033
rect 18843 44347 18909 44963
rect 19365 45027 19435 45033
rect 19365 44642 19435 44959
rect 19941 44784 20003 45025
rect 19936 44779 20008 44784
rect 19936 44723 19941 44779
rect 20003 44723 20008 44779
rect 19936 44718 20008 44723
rect 19360 44637 19440 44642
rect 19360 44567 19365 44637
rect 19435 44567 19440 44637
rect 19360 44562 19440 44567
rect 18838 44342 18914 44347
rect 18838 44286 18843 44342
rect 18909 44286 18914 44342
rect 18838 44281 18914 44286
rect 1636 44149 1702 44151
rect 1531 44148 1707 44149
rect 1354 44146 1707 44148
rect 1354 44090 1641 44146
rect 1697 44090 1707 44146
rect 1354 44088 1707 44090
rect 396 43994 402 44058
rect 466 44056 472 44058
rect 1354 44056 1414 44088
rect 1531 44087 1707 44088
rect 1636 44085 1702 44087
rect 466 43996 1414 44056
rect 466 43994 472 43996
rect 950 43569 956 43633
rect 1020 43631 1026 43633
rect 4258 43631 4324 43634
rect 1020 43629 4324 43631
rect 1020 43573 4263 43629
rect 4319 43573 4324 43629
rect 1020 43571 4324 43573
rect 1020 43569 1026 43571
rect 4258 43568 4324 43571
<< via3 >>
rect 18843 44963 18909 45027
rect 19365 44959 19435 45027
rect 402 43994 466 44058
rect 956 43569 1020 43633
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 45028 18890 45152
rect 19382 45028 19442 45152
rect 18830 45027 18910 45028
rect 18830 44963 18843 45027
rect 18909 44963 18910 45027
rect 18830 44962 18910 44963
rect 19364 45027 19442 45028
rect 18830 44952 18890 44962
rect 19364 44959 19365 45027
rect 19435 44959 19442 45027
rect 19364 44958 19442 44959
rect 19382 44952 19442 44958
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 44058 600 44152
rect 200 43994 402 44058
rect 466 43994 600 44058
rect 200 1000 600 43994
rect 800 43633 1200 44152
rect 800 43569 956 43633
rect 1020 43569 1200 43633
rect 800 1000 1200 43569
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use manchester_decoder  manchester_decoder_0
timestamp 1738528573
transform 1 0 6086 0 1 43632
box -38 -48 682 592
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1200 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22634 0 22814 200 0 FreeSans 1200 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18770 0 18950 200 0 FreeSans 1200 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 14906 0 15086 200 0 FreeSans 1200 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 11042 0 11222 200 0 FreeSans 1200 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 7178 0 7358 200 0 FreeSans 1200 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 3314 0 3494 200 0 FreeSans 1200 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 200 1000 600 44152 1 FreeSans 500 0 0 0 VDPWR
port 52 nsew
flabel metal4 s 800 1000 1200 44152 1 FreeSans 500 0 0 0 VGND
port 53 nsew
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 34 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
