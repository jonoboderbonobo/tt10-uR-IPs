magic
tech sky130A
magscale 1 2
timestamp 1741560675
<< nwell >>
rect 598 1140 634 1246
rect 1154 1140 1188 1246
rect 1701 1140 2038 1246
rect 66 970 2254 1140
rect 598 794 634 970
rect 1154 794 1188 970
rect 598 713 1493 794
rect 603 700 1493 713
rect 605 699 890 700
rect 1160 699 1424 700
rect 1701 699 2038 970
<< poly >>
rect -18 688 48 698
rect -18 654 -2 688
rect 32 654 96 688
rect 564 654 665 688
rect 1126 654 1220 688
rect 1670 654 1775 688
rect -18 644 48 654
<< polycont >>
rect -2 654 32 688
<< locali >>
rect -2 688 32 704
rect -2 638 32 654
rect 445 17 2188 51
<< viali >>
rect -2 654 32 688
<< metal1 >>
rect -20 1228 2174 1261
rect -20 1227 1064 1228
rect 443 1222 1064 1227
rect 459 1210 497 1222
rect 1014 1210 1064 1222
rect 1052 1201 1064 1210
rect 1553 1201 1619 1228
rect 2108 1202 2174 1228
rect 498 1054 550 1060
rect 498 996 550 1002
rect 1058 1054 1110 1060
rect 1058 996 1110 1002
rect 1615 1054 1667 1060
rect 2155 1002 2161 1054
rect 2213 1002 2219 1054
rect 1615 996 1667 1002
rect -20 688 38 704
rect -20 654 -2 688
rect 32 654 38 688
rect -20 638 38 654
rect 572 648 631 695
rect 1131 694 1186 695
rect 1128 648 1186 694
rect 1666 648 1741 695
rect 485 311 491 363
rect 543 311 549 363
rect -20 51 80 52
rect -20 16 447 51
rect 603 1 631 648
rect 1040 363 1092 369
rect 1040 305 1092 311
rect 1158 1 1186 648
rect 1615 363 1667 369
rect 1615 305 1667 311
rect 1713 1 1741 648
rect 2171 363 2223 369
rect 2171 305 2223 311
<< via1 >>
rect 498 1002 550 1054
rect 1058 1002 1110 1054
rect 1615 1002 1667 1054
rect 2161 1002 2213 1054
rect 491 311 543 363
rect 1040 311 1092 363
rect 1615 311 1667 363
rect 2171 311 2223 363
<< metal2 >>
rect 2161 1054 2213 1060
rect 492 1042 498 1054
rect -20 1014 498 1042
rect 492 1002 498 1014
rect 550 1042 556 1054
rect 1052 1042 1058 1054
rect 550 1014 1058 1042
rect 550 1002 556 1014
rect 1052 1002 1058 1014
rect 1110 1042 1116 1054
rect 1609 1042 1615 1054
rect 1110 1014 1615 1042
rect 1110 1002 1116 1014
rect 1609 1002 1615 1014
rect 1667 1042 1673 1054
rect 1667 1014 2161 1042
rect 1667 1002 1673 1014
rect 2161 996 2213 1002
rect 491 363 543 369
rect -20 323 491 351
rect 1034 351 1040 363
rect 543 323 1040 351
rect 1034 311 1040 323
rect 1092 351 1098 363
rect 1609 351 1615 363
rect 1092 323 1615 351
rect 1092 311 1098 323
rect 1609 311 1615 323
rect 1667 351 1673 363
rect 2165 351 2171 363
rect 1667 323 2171 351
rect 1667 311 1673 323
rect 2165 311 2171 323
rect 2223 311 2229 363
rect 491 305 543 311
use schmTrigg  stage_1 schmTrig
timestamp 1741560675
transform 1 0 793 0 1 2064
box 934 -2152 1557 -803
use schmTrigg  stage_2
timestamp 1741560675
transform 1 0 -872 0 1 2064
box 934 -2152 1557 -803
use schmTrigg  stage_3
timestamp 1741560675
transform 1 0 -317 0 1 2064
box 934 -2152 1557 -803
use schmTrigg  stage_out
timestamp 1741560675
transform 1 0 238 0 1 2064
box 934 -2152 1557 -803
<< end >>
