** sch_path: /foss/designs/tt10-uR-IPs/xschem/breakdown_voltage_tb.sch
**.subckt breakdown_voltage_tb
.save v(in)
.save v(out)
XM2 in in out GND sky130_fd_pr__nfet_01v8 L=0.15 W=30 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
Vdrain in GND 3
XR10 GND out GND sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
**** begin user architecture code


.control
*set filetype=ascii
*save all

op
DC Vdrain 0 500 1


write tb_breakdown_voltage.raw
*exit

.endc



** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
