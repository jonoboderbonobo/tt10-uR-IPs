magic
tech sky130A
magscale 1 2
timestamp 1741560675
<< nwell >>
rect 24539 3976 24722 3978
<< locali >>
rect 25887 3741 25921 4056
<< viali >>
rect 25887 3707 25921 3741
<< metal1 >>
rect 25757 4832 25785 5198
rect 24640 4804 25785 4832
rect 24640 4643 24668 4804
rect 27984 4585 28567 4633
rect 24277 4460 24341 4466
rect 24277 4408 24283 4460
rect 24335 4448 24341 4460
rect 24335 4420 24597 4448
rect 24335 4408 24341 4420
rect 24277 4402 24341 4408
rect 25168 4302 25220 4308
rect 25168 4244 25220 4250
rect 25767 3997 25819 4003
rect 25767 3939 25819 3945
rect 26371 3997 26423 4003
rect 26371 3939 26423 3945
rect 26926 3997 26978 4003
rect 26926 3939 26978 3945
rect 27481 3997 27533 4003
rect 27481 3939 27533 3945
rect 26938 3938 26966 3939
rect 28519 3796 28567 4585
rect 28519 3750 28568 3796
rect 25875 3741 25933 3747
rect 25875 3707 25887 3741
rect 25921 3707 25933 3741
rect 25875 3701 25933 3707
rect 25887 1483 25921 3701
rect 25887 1449 26621 1483
rect 26587 1038 26621 1449
rect 28520 1482 28568 3750
rect 28520 1434 30442 1482
rect 26498 894 26678 1038
rect 30394 984 30442 1434
rect 26492 714 26498 894
rect 26678 714 26684 894
rect 30362 732 30542 984
rect 30356 552 30362 732
rect 30542 552 30548 732
<< via1 >>
rect 24283 4408 24335 4460
rect 25168 4250 25220 4302
rect 25767 3945 25819 3997
rect 26371 3945 26423 3997
rect 26926 3945 26978 3997
rect 27481 3945 27533 3997
rect 26498 714 26678 894
rect 30362 552 30542 732
<< metal2 >>
rect 24217 4951 25791 4979
rect 24217 4471 24245 4951
rect 25116 4491 25296 4519
rect 24203 4466 24277 4471
rect 24203 4462 24341 4466
rect 24203 4406 24212 4462
rect 24268 4460 24341 4462
rect 24268 4408 24283 4460
rect 24335 4408 24341 4460
rect 24268 4406 24341 4408
rect 24203 4402 24341 4406
rect 24203 4397 24277 4402
rect 25053 4246 25062 4302
rect 25118 4288 25127 4302
rect 25162 4288 25168 4302
rect 25118 4260 25168 4288
rect 25118 4246 25127 4260
rect 25162 4250 25168 4260
rect 25220 4250 25226 4302
rect 25268 3985 25296 4491
rect 25324 4246 25333 4302
rect 25389 4288 25398 4302
rect 25389 4260 25785 4288
rect 25389 4246 25398 4260
rect 25761 3985 25767 3997
rect 25268 3957 25767 3985
rect 25761 3945 25767 3957
rect 25819 3945 25825 3997
rect 26365 3945 26371 3997
rect 26423 3945 26429 3997
rect 26920 3945 26926 3997
rect 26978 3945 26984 3997
rect 27475 3945 27481 3997
rect 27533 3988 27539 3997
rect 27533 3954 27762 3988
rect 27533 3945 27539 3954
rect 26383 3762 26411 3945
rect 26920 3939 26984 3945
rect 26938 3762 26966 3939
rect 27734 3762 27762 3954
rect 26360 3706 26369 3762
rect 26425 3706 26434 3762
rect 26915 3706 26924 3762
rect 26980 3706 26989 3762
rect 27711 3706 27720 3762
rect 27776 3706 27785 3762
rect 26498 894 26678 900
rect 26498 527 26678 714
rect 30362 732 30542 738
rect 26494 357 26503 527
rect 26673 357 26682 527
rect 30362 519 30542 552
rect 26498 352 26678 357
rect 30358 349 30367 519
rect 30537 349 30546 519
rect 30362 344 30542 349
<< via2 >>
rect 24212 4406 24268 4462
rect 25062 4246 25118 4302
rect 25333 4246 25389 4302
rect 26369 3706 26425 3762
rect 26924 3706 26980 3762
rect 27720 3706 27776 3762
rect 26503 357 26673 527
rect 30367 349 30537 519
<< metal3 >>
rect 410 4466 486 4472
rect 410 4402 416 4466
rect 480 4464 486 4466
rect 24203 4464 24273 4467
rect 480 4462 24273 4464
rect 480 4406 24212 4462
rect 24268 4406 24273 4462
rect 480 4404 24273 4406
rect 480 4402 486 4404
rect 410 4396 486 4402
rect 24203 4401 24273 4404
rect 24134 4242 24140 4306
rect 24204 4304 24210 4306
rect 25057 4304 25123 4307
rect 25328 4304 25394 4307
rect 24204 4302 25394 4304
rect 24204 4246 25062 4302
rect 25118 4246 25333 4302
rect 25389 4246 25394 4302
rect 24204 4244 25394 4246
rect 24204 4242 24210 4244
rect 25057 4241 25123 4244
rect 25328 4241 25394 4244
rect 26367 3767 26427 4076
rect 26692 4017 26982 4067
rect 26922 3767 26982 4017
rect 27718 3767 27778 4091
rect 26364 3762 26430 3767
rect 26364 3706 26369 3762
rect 26425 3706 26430 3762
rect 26364 3701 26430 3706
rect 26919 3762 26985 3767
rect 26919 3706 26924 3762
rect 26980 3706 26985 3762
rect 26919 3701 26985 3706
rect 27715 3762 27781 3767
rect 27715 3706 27720 3762
rect 27776 3706 27781 3762
rect 27715 3701 27781 3706
rect 26498 527 26678 532
rect 26498 357 26503 527
rect 26673 357 26678 527
rect 26498 213 26678 357
rect 26498 172 26562 213
rect 26556 149 26562 172
rect 26626 172 26678 213
rect 30362 519 30542 524
rect 30362 349 30367 519
rect 30537 349 30542 519
rect 30362 220 30542 349
rect 30362 198 30410 220
rect 26626 149 26632 172
rect 30404 156 30410 198
rect 30474 198 30542 220
rect 30474 156 30480 198
rect 30404 150 30480 156
rect 26556 143 26632 149
<< via3 >>
rect 416 4402 480 4466
rect 24140 4242 24204 4306
rect 26562 149 26626 213
rect 30410 156 30474 220
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 4466 600 44152
rect 200 4402 416 4466
rect 480 4402 600 4466
rect 200 1000 600 4402
rect 800 4304 1200 44152
rect 24139 4997 28127 5057
rect 24139 4996 25826 4997
rect 24139 4307 24200 4996
rect 24139 4306 24205 4307
rect 24139 4304 24140 4306
rect 800 4244 24140 4304
rect 800 1000 1200 4244
rect 24139 4242 24140 4244
rect 24204 4242 24205 4306
rect 24139 4241 24205 4242
rect 30404 220 30480 226
rect 26556 213 26632 219
rect 26556 200 26562 213
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 149 26562 200
rect 26626 200 26632 213
rect 30404 200 30410 220
rect 26626 149 26678 200
rect 26498 0 26678 149
rect 30362 156 30410 200
rect 30474 200 30480 220
rect 30474 156 30542 200
rect 30362 0 30542 156
use ibias_10nA  bias /foss/designs/tt10-uR-IPs/magic/tt10/biasGen
timestamp 1741558662
transform 1 0 24418 0 1 5576
box 5 -1612 850 -838
use s130_mim_sl_40fF  cap_osc_1 /foss/designs/tt10-uR-IPs/magic/tt10/osc/cap
timestamp 1741556153
transform 1 0 28037 0 1 4636
box -474 -628 182 628
use s130_mim_sl_40fF  cap_osc_2
timestamp 1741556153
transform 1 0 26230 0 1 4636
box -474 -628 182 628
use s130_mim_sl_40fF  cap_osc_3
timestamp 1741556153
transform 1 0 27141 0 1 4646
box -474 -628 182 628
use osc  osc_0 /foss/designs/tt10-uR-IPs/magic/tt10/osc
timestamp 1741560675
transform 1 0 25777 0 1 3937
box -20 -88 2350 1261
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
