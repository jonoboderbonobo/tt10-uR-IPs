** sch_path: /foss/designs/tt10-uR-IPs/xschem/T2/biasGen/A_tt10_10nA/ibias_10nA_PARAX_tran_tb.sch
**.subckt ibias_10nA_PARAX_tran_tb
VIN1 net1 0 0 pulse 0 1.8 10m 1m 1m 10m 20m ac 1 0
vi_total net1 VDD_jump 0
.save i(vi_total)
vi_d V1 net2 0
.save i(vi_d)
x1 VDD_jump 0 Vnbias Vpbias ibias_10nA
XM55 V1 Vpbias VDD_jump VDD_jump sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R25 net2 V3 10k m=1
XM2 V3 Vnbias V4 V4 sky130_fd_pr__nfet_01v8 L=0.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
vi_d1 V4 0 0
.save i(vi_d1)
vi_d_parax V1_parax net3 0
.save i(vi_d_parax)
XM1 V1_parax Vpbias_parax VDD_jump VDD_jump sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R24 net3 V3_parax 10k m=1
XM3 V3_parax Vnbias_parax V4_parax V4_parax sky130_fd_pr__nfet_01v8 L=0.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
vi_d3 V4_parax 0 0
.save i(vi_d3)
x2 VDD_jump 0 Vnbias_parax Vpbias_parax ibias_10nA_parax
**** begin user architecture code



.temp 30

*.option gmin=5n
*.option scale=1e-6
.option wnflag=1
.option savecurrents

.save all
.control
  save all alli
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm1.msky130_fd_pr__nfet_01v8[id]
  save @m.xm1.msky130_fd_pr__nfet_01v8[vgs]

  save @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
  save @m.xm1.msky130_fd_pr__nfet_01v8[cgs]
  save @m.xm1.msky130_fd_pr__nfet_01v8[cgdo]
  save @m.xm1.msky130_fd_pr__nfet_01v8[cgb]

  save @m.xm1.msky130_fd_pr__nfet_01v8[vds]
  save @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
  save @m.xm1.msky130_fd_pr__nfet_01v8[vth]


  save @m.xm1.msky130_fd_pr__nfet_01v8[leff]
  save @m.xm1.msky130_fd_pr__nfet_01v8[weff]
  save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
  save @m.xm1.msky130_fd_pr__nfet_01v8[l]
  save @m.xm1.msky130_fd_pr__nfet_01v8[w]
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]








  tran 1m 50m
  remzerovec
  write nmos_tb_tran.raw

  op
  set appendwrite
  remzerovec
  write nmos_tb_tran.raw






  *quit 0




.endc




** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


**** end user architecture code
**.ends

* expanding   symbol:  T2/biasGen/A_tt10_10nA/ibias_10nA.sym # of pins=4
** sym_path: /foss/designs/tt10-uR-IPs/xschem/T2/biasGen/A_tt10_10nA/ibias_10nA.sym
** sch_path: /foss/designs/tt10-uR-IPs/xschem/T2/biasGen/A_tt10_10nA/ibias_10nA.sch
.subckt ibias_10nA Vdd Vss Vnbias Vpbias
*.ipin Vdd
*.ipin Vss
*.opin Vnbias
*.opin Vpbias
XM3 Vpbias Vpbias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vnbias Vpbias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 Vpbias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vpbias Vnbias net1 Vss sky130_fd_pr__nfet_01v8 L=0.2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vnbias Vnbias Vss Vss sky130_fd_pr__nfet_01v8 L=0.2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 net2 net1 Vss sky130_fd_pr__nfet_01v8 L=0.2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net1 net2 Vss Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  T2/biasGen/A_tt10_10nA/ibias_10nA_parax.sym # of pins=4
** sym_path: /foss/designs/tt10-uR-IPs/xschem/T2/biasGen/A_tt10_10nA/ibias_10nA_parax.sym
.include T2/biasGen/A_tt10_10nA/ibias_10nA_parax.spice
.end
