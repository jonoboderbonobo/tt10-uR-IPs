magic
tech sky130A
magscale 1 2
timestamp 1738157446
<< checkpaint >>
rect -86 -651 2856 -598
rect -86 -704 3225 -651
rect -86 -3938 3594 -704
rect 283 -3991 3594 -3938
rect 652 -4044 3594 -3991
<< error_s >>
rect 338 -951 373 -917
rect 339 -970 373 -951
rect 191 -1200 200 -1072
rect 219 -1228 228 -1100
rect 147 -2347 209 -2341
rect 147 -2381 159 -2347
rect 147 -2387 209 -2381
rect 358 -2483 373 -970
rect 392 -1004 427 -970
rect 747 -1004 782 -970
rect 392 -2483 426 -1004
rect 748 -1023 782 -1004
rect 556 -1072 618 -1066
rect 556 -1106 568 -1072
rect 556 -1112 618 -1106
rect 556 -2400 618 -2394
rect 556 -2434 568 -2400
rect 556 -2440 618 -2434
rect 392 -2517 407 -2483
rect 767 -2536 782 -1023
rect 801 -1057 836 -1023
rect 801 -2536 835 -1057
rect 965 -1125 1027 -1119
rect 965 -1159 977 -1125
rect 965 -1165 1027 -1159
rect 1157 -1858 1191 -1840
rect 1157 -1894 1227 -1858
rect 1174 -1928 1245 -1894
rect 1525 -1928 1560 -1894
rect 965 -2453 1027 -2447
rect 965 -2487 977 -2453
rect 965 -2493 1027 -2487
rect 801 -2570 816 -2536
rect 1174 -2589 1244 -1928
rect 1526 -1947 1560 -1928
rect 1356 -1996 1414 -1990
rect 1356 -2030 1368 -1996
rect 1356 -2036 1414 -2030
rect 1356 -2506 1414 -2500
rect 1356 -2540 1368 -2506
rect 1356 -2546 1414 -2540
rect 1174 -2625 1227 -2589
rect 1545 -2642 1560 -1947
rect 1579 -1981 1614 -1947
rect 1579 -2642 1613 -1981
rect 1725 -2049 1783 -2043
rect 1725 -2083 1737 -2049
rect 1725 -2089 1783 -2083
rect 1725 -2559 1783 -2553
rect 1725 -2593 1737 -2559
rect 1725 -2599 1783 -2593
rect 1579 -2676 1594 -2642
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_lvt_3YHUUE  XM1
timestamp 0
transform 1 0 1754 0 1 -2321
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_2NKB8S  XM2
timestamp 0
transform 1 0 587 0 1 -1753
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_3YHUUE  XM3
timestamp 0
transform 1 0 2123 0 1 -2374
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_2NKB8S  XM4
timestamp 0
transform 1 0 996 0 1 -1806
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_3YHUUE  XM6
timestamp 0
transform 1 0 1385 0 1 -2268
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_2NKB8S  XM10
timestamp 0
transform 1 0 178 0 1 -1700
box -231 -819 231 819
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vss
port 3 nsew
<< end >>
