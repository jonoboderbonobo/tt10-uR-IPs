** sch_path: /tmp/xschem_web_dcfaafabed/BGR_SKY130_final.sch
**.subckt BGR_SKY130_final
XM1 net2 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S1*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 net8 net2 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S2*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net7 net8 net1 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S3*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net4 net5 net1 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S4*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net5 net5 net4 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S5*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net3 net6 net4 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S6*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net6 net6 net3 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S7*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net7 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S8*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net8 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S9*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net5 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S10*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net6 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S11*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net9 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S12*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMc net10 net11 net3 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S15*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMb net11 net11 net10 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S14*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMa net11 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S13*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMf net9 net12 net10 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S18*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMe net12 net12 net9 GND sky130_fd_pr__nfet_01v8_lvt L={L} W={S17*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMd net12 net7 VDD VDD sky130_fd_pr__pfet_01v8_lvt L={L} W={S16*L} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 VDD GND 1.8
C1 net9 GND 1p m=1
XQ1 GND GND net8 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
**** begin user architecture code


** Analysis Requests **
.op
** Outputs Requests **
.control
run
show > opota.txt
.endc


 ** manual skywater pdks install (with patches applied)
*.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0

.include /foss/pdks/sky130A/libs.tech/combined/sky130_fd_pr__model__pnp.model.spice



** Analysis Requests **
** Outputs Requests **
.control
dc temp -40 125 5 V1 1.2 2.2 0.1
plot V(net2)
plot V(net8)

plot V(net9)
.endc




.param L = 1

*** 1st Branch: Controls amount of current in Bjt
.param S9 = 15

*** 2nd Branch:Controls Initial Offset
.param S8 = 1
.param S3 = 64
.param S2 = 64
.param S1 = 64

*** 3rd, 4th, 5th Branches: Fine Tuning slope for PTAT slope
.param S10 = 1
.param S5 = 4
.param S4 = 1

.param S11 = 1
.param S7 = 4
.param S6 = 1


.param S13 = 1
.param S14 = 4
.param S15 = 1

.param S16 = 1
.param S17 = 4
.param S18 = 1

*** Branch 6: Coarse Tuning for PTAT Slope
.param S12 = 1


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
