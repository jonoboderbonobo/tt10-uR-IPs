magic
tech sky130A
magscale 1 2
timestamp 1741523581
<< locali >>
rect 27845 1407 27879 1722
<< viali >>
rect 27845 1373 27879 1407
<< metal1 >>
rect 27381 2830 27758 2864
rect 26470 2344 26476 2396
rect 26528 2344 26534 2396
rect 26932 2145 26938 2197
rect 26990 2145 26996 2197
rect 26364 2047 26370 2099
rect 26422 2096 26428 2099
rect 26422 2050 26512 2096
rect 26422 2047 26428 2050
rect 26476 1533 26522 1667
rect 27381 1533 27427 2830
rect 29942 2251 30525 2299
rect 27705 1659 27757 1665
rect 27705 1601 27757 1607
rect 28338 1590 28366 1632
rect 28893 1598 28921 1632
rect 29448 1602 29476 1632
rect 28881 1592 28933 1598
rect 26476 1487 27427 1533
rect 28326 1584 28378 1590
rect 28881 1534 28933 1540
rect 29436 1596 29488 1602
rect 29436 1538 29488 1544
rect 28326 1526 28378 1532
rect 27833 1407 27891 1413
rect 27833 1373 27845 1407
rect 27879 1373 27891 1407
rect 27833 1367 27891 1373
rect 26498 1077 26678 1106
rect 27845 1077 27879 1367
rect 26498 1043 27879 1077
rect 26498 894 26678 1043
rect 30477 984 30525 2251
rect 26492 714 26498 894
rect 26678 714 26684 894
rect 30362 732 30542 984
rect 30356 552 30362 732
rect 30542 552 30548 732
<< via1 >>
rect 26476 2344 26528 2396
rect 26938 2145 26990 2197
rect 26370 2047 26422 2099
rect 27705 1607 27757 1659
rect 28326 1532 28378 1584
rect 28881 1540 28933 1592
rect 29436 1544 29488 1596
rect 26498 714 26678 894
rect 30362 552 30542 732
<< metal2 >>
rect 26175 2617 27749 2645
rect 26175 2133 26203 2617
rect 26372 2343 26381 2399
rect 26437 2386 26446 2399
rect 26476 2396 26528 2402
rect 26437 2355 26476 2386
rect 26437 2343 26446 2355
rect 26476 2338 26528 2344
rect 26938 2197 26990 2203
rect 26990 2148 27321 2194
rect 26938 2139 26990 2145
rect 26175 2128 26221 2133
rect 26161 2072 26170 2128
rect 26226 2096 26235 2128
rect 26370 2099 26422 2105
rect 26226 2072 26370 2096
rect 26175 2050 26370 2072
rect 26370 2041 26422 2047
rect 27275 1656 27321 2148
rect 27449 1912 27458 1968
rect 27514 1954 27523 1968
rect 27514 1926 27743 1954
rect 27514 1912 27523 1926
rect 27699 1656 27705 1659
rect 27275 1610 27705 1656
rect 27699 1607 27705 1610
rect 27757 1607 27763 1659
rect 28320 1532 28326 1584
rect 28378 1532 28384 1584
rect 28875 1540 28881 1592
rect 28933 1540 28939 1592
rect 29430 1544 29436 1596
rect 29488 1544 29494 1596
rect 28338 1441 28366 1532
rect 28324 1432 28380 1441
rect 28893 1439 28921 1540
rect 28324 1367 28380 1376
rect 28879 1430 28935 1439
rect 29448 1423 29476 1544
rect 28879 1365 28935 1374
rect 29434 1414 29490 1423
rect 29434 1349 29490 1358
rect 26498 894 26678 900
rect 26498 527 26678 714
rect 30362 732 30542 738
rect 26494 357 26503 527
rect 26673 357 26682 527
rect 30362 519 30542 552
rect 26498 352 26678 357
rect 30358 349 30367 519
rect 30537 349 30546 519
rect 30362 344 30542 349
<< via2 >>
rect 26381 2343 26437 2399
rect 26170 2072 26226 2128
rect 27458 1912 27514 1968
rect 28324 1376 28380 1432
rect 28879 1374 28935 1430
rect 29434 1358 29490 1414
rect 26503 357 26673 527
rect 30367 349 30537 519
<< metal3 >>
rect 26376 2401 26442 2404
rect 25850 2399 26442 2401
rect 25850 2343 26381 2399
rect 26437 2343 26442 2399
rect 25850 2341 26442 2343
rect 25408 2129 25472 2135
rect 370 2065 376 2129
rect 440 2127 446 2129
rect 440 2067 25408 2127
rect 440 2065 446 2067
rect 25408 2059 25472 2065
rect 25850 2034 25910 2341
rect 26376 2338 26442 2341
rect 26002 2068 26008 2132
rect 26072 2130 26078 2132
rect 26165 2130 26231 2133
rect 26072 2128 26231 2130
rect 26072 2072 26170 2128
rect 26226 2072 26231 2128
rect 26072 2070 26231 2072
rect 26072 2068 26078 2070
rect 26165 2067 26231 2070
rect 25760 1970 25766 1972
rect 25752 1910 25766 1970
rect 25760 1908 25766 1910
rect 25830 1970 25910 2034
rect 27453 1970 27519 1973
rect 25830 1968 27519 1970
rect 25830 1912 27458 1968
rect 27514 1912 27519 1968
rect 25830 1910 27519 1912
rect 25830 1908 25836 1910
rect 27453 1907 27519 1910
rect 28319 1434 28385 1437
rect 28502 1434 28562 1788
rect 28319 1432 28562 1434
rect 28319 1376 28324 1432
rect 28380 1376 28562 1432
rect 28319 1374 28562 1376
rect 28874 1432 28940 1435
rect 29164 1432 29224 1796
rect 28874 1430 29224 1432
rect 28874 1374 28879 1430
rect 28935 1374 29224 1430
rect 28319 1371 28385 1374
rect 28874 1372 29224 1374
rect 29429 1416 29495 1419
rect 30630 1416 30690 1786
rect 29429 1414 30690 1416
rect 28874 1369 28940 1372
rect 29429 1358 29434 1414
rect 29490 1358 30690 1414
rect 29429 1356 30690 1358
rect 29429 1353 29495 1356
rect 26498 527 26678 532
rect 26498 357 26503 527
rect 26673 357 26678 527
rect 26498 199 26678 357
rect 30362 519 30542 524
rect 30362 349 30367 519
rect 30537 349 30542 519
rect 30362 199 30542 349
rect 26493 21 26499 199
rect 26677 21 26683 199
rect 30357 21 30363 199
rect 30541 21 30547 199
rect 26498 20 26678 21
rect 30362 20 30542 21
<< via3 >>
rect 376 2065 440 2129
rect 25408 2065 25472 2129
rect 26008 2068 26072 2132
rect 25766 1908 25830 1972
rect 26499 21 26677 199
rect 30363 21 30541 199
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 2129 600 44152
rect 200 2065 376 2129
rect 440 2065 600 2129
rect 200 1000 600 2065
rect 800 1970 1200 44152
rect 24193 2953 30549 3015
rect 24193 1970 24255 2953
rect 26002 2132 26073 2133
rect 25407 2129 25473 2130
rect 25407 2065 25408 2129
rect 25472 2127 25473 2129
rect 26002 2127 26008 2132
rect 25472 2068 26008 2127
rect 26072 2068 26073 2132
rect 25472 2067 26073 2068
rect 25472 2065 25473 2067
rect 25407 2064 25473 2065
rect 25765 1972 25831 1973
rect 25765 1970 25766 1972
rect 800 1910 25766 1970
rect 800 1000 1200 1910
rect 25765 1908 25766 1910
rect 25830 1908 25831 1972
rect 25765 1907 25831 1908
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 199 26678 200
rect 26498 21 26499 199
rect 26677 21 26678 199
rect 26498 0 26678 21
rect 30362 199 30542 200
rect 30362 21 30363 199
rect 30541 21 30542 199
rect 30362 0 30542 21
use ibias_10nA  ibias_10nA_0 /foss/designs/tt10-uR-IPs/magic/tt10/biasGen
timestamp 1741378290
transform 1 0 26376 0 1 3242
box -92 -1634 850 -857
use osc  osc_0 /foss/designs/tt10-uR-IPs/magic/tt10/osc
timestamp 1741465372
transform 1 0 27735 0 1 1603
box -20 1 2272 1261
use sky130_fd_pr__cap_mim_m3_1_2BN6ET  sky130_fd_pr__cap_mim_m3_1_2BN6ET_0
timestamp 1741467963
transform 0 -1 29598 1 0 2354
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_2BN6ET  sky130_fd_pr__cap_mim_m3_1_2BN6ET_1
timestamp 1741467963
transform 0 -1 28290 1 0 2354
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_2BN6ET  sky130_fd_pr__cap_mim_m3_1_2BN6ET_2
timestamp 1741467963
transform 0 -1 30908 1 0 2354
box -686 -540 686 540
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
