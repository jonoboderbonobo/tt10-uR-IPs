magic
tech sky130A
magscale 1 2
timestamp 1738518703
<< viali >>
rect 6288 43847 6322 43881
rect 6515 43847 6549 43881
rect 6661 43726 6695 43760
<< metal1 >>
rect 6086 44223 6117 44224
rect 5815 44221 6117 44223
rect 1984 44196 6117 44221
rect 1984 44194 6088 44196
rect 1984 44193 6030 44194
rect 1787 44091 1793 44143
rect 1845 44133 1851 44143
rect 1984 44133 2012 44193
rect 5815 44192 6030 44193
rect 1845 44100 2015 44133
rect 1845 44091 1851 44100
rect 5795 43896 5857 43902
rect 7027 43900 7097 43906
rect 5857 43881 6338 43896
rect 5857 43847 6288 43881
rect 6322 43847 6338 43881
rect 5857 43836 6338 43847
rect 6500 43881 7027 43900
rect 6500 43847 6515 43881
rect 6549 43847 7027 43881
rect 5857 43834 6300 43836
rect 5795 43828 5857 43834
rect 6500 43830 7027 43847
rect 7027 43824 7097 43830
rect 6642 43779 6800 43780
rect 7271 43779 7337 43785
rect 6642 43760 7271 43779
rect 6642 43726 6661 43760
rect 6695 43726 7271 43760
rect 6642 43713 7271 43726
rect 6642 43712 6800 43713
rect 7271 43707 7337 43713
rect 4463 43574 4469 43626
rect 4521 43615 4527 43626
rect 4521 43584 6126 43615
rect 4521 43574 4527 43584
<< via1 >>
rect 1793 44091 1845 44143
rect 5795 43834 5857 43896
rect 7027 43830 7097 43900
rect 7271 43713 7337 43779
rect 4469 43574 4521 43626
<< metal2 >>
rect 7027 44771 7097 44780
rect 5792 44703 5801 44765
rect 5857 44703 5866 44765
rect 1632 44090 1641 44146
rect 1697 44134 1706 44146
rect 1793 44143 1845 44149
rect 1697 44101 1793 44134
rect 1697 44090 1706 44101
rect 1793 44085 1845 44091
rect 5795 43896 5857 44703
rect 7027 43900 7097 44711
rect 7271 44453 7337 44462
rect 5789 43834 5795 43896
rect 5857 43834 5863 43896
rect 7021 43830 7027 43900
rect 7097 43830 7103 43900
rect 7271 43779 7337 44397
rect 7265 43713 7271 43779
rect 7337 43713 7343 43779
rect 4263 43629 4319 43638
rect 4469 43626 4521 43632
rect 4319 43585 4469 43616
rect 4263 43564 4319 43573
rect 4469 43568 4521 43574
<< via2 >>
rect 5801 44703 5857 44765
rect 7027 44711 7097 44771
rect 1641 44090 1697 44146
rect 7271 44397 7337 44453
rect 4263 43573 4319 43629
<< metal3 >>
rect 7227 45041 7293 45047
rect 6685 45025 6755 45031
rect 6132 45012 6196 45018
rect 6132 44942 6196 44948
rect 5796 44765 5862 44770
rect 6133 44765 6195 44942
rect 5796 44703 5801 44765
rect 5857 44703 6195 44765
rect 6685 44776 6755 44957
rect 6685 44771 7102 44776
rect 6685 44711 7027 44771
rect 7097 44711 7102 44771
rect 6685 44706 7102 44711
rect 5796 44698 5862 44703
rect 7227 44458 7293 44977
rect 7227 44453 7342 44458
rect 7227 44397 7271 44453
rect 7337 44397 7342 44453
rect 7227 44392 7342 44397
rect 1636 44149 1702 44151
rect 1531 44148 1707 44149
rect 1354 44146 1707 44148
rect 1354 44090 1641 44146
rect 1697 44090 1707 44146
rect 1354 44088 1707 44090
rect 396 43994 402 44058
rect 466 44056 472 44058
rect 1354 44056 1414 44088
rect 1531 44087 1707 44088
rect 1636 44085 1702 44087
rect 466 43996 1414 44056
rect 466 43994 472 43996
rect 950 43569 956 43633
rect 1020 43631 1026 43633
rect 4258 43631 4324 43634
rect 1020 43629 4324 43631
rect 1020 43573 4263 43629
rect 4319 43573 4324 43629
rect 1020 43571 4324 43573
rect 1020 43569 1026 43571
rect 4258 43568 4324 43571
<< via3 >>
rect 6132 44948 6196 45012
rect 6685 44957 6755 45025
rect 7227 44977 7293 45041
rect 402 43994 466 44058
rect 956 43569 1020 43633
<< metal4 >>
rect 6134 45013 6194 45152
rect 6686 45026 6746 45152
rect 7238 45042 7298 45152
rect 7226 45041 7298 45042
rect 6684 45025 6756 45026
rect 6131 45012 6197 45013
rect 6131 44948 6132 45012
rect 6196 44948 6197 45012
rect 6684 44957 6685 45025
rect 6755 44957 6756 45025
rect 7226 44977 7227 45041
rect 7293 44977 7298 45041
rect 7226 44976 7298 44977
rect 6684 44956 6756 44957
rect 6686 44952 6746 44956
rect 7238 44952 7298 44976
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 6131 44947 6197 44948
rect 200 44058 600 44152
rect 200 43994 402 44058
rect 466 43994 600 44058
rect 200 1000 600 43994
rect 800 43633 1200 44152
rect 800 43569 956 43633
rect 1020 43569 1200 43633
rect 800 1000 1200 43569
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use manchester_decoder  manchester_decoder_0
timestamp 1738500547
transform 1 0 6086 0 1 43632
box -38 -48 682 592
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
