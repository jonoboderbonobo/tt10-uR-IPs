magic
tech sky130A
magscale 1 2
timestamp 1741541561
<< nwell >>
rect 934 -842 1479 -818
rect 934 -847 1234 -842
rect 1143 -851 1234 -847
rect 1152 -894 1234 -851
rect 1315 -847 1479 -842
rect 1152 -895 1291 -894
rect 1315 -895 1453 -847
rect 1152 -997 1453 -895
rect 1064 -1056 1104 -1050
rect 1064 -1077 1110 -1056
rect 1145 -1072 1453 -997
rect 1145 -1074 1239 -1072
rect 1145 -1082 1223 -1074
rect 1284 -1180 1453 -1072
rect 1284 -1184 1464 -1180
rect 1230 -1195 1464 -1184
rect 1230 -1365 1479 -1195
<< poly >>
rect 1028 -1129 1058 -1075
rect 1028 -1376 1058 -1329
rect 1115 -1359 1145 -1329
rect 934 -1410 1058 -1376
rect 1028 -1422 1058 -1410
rect 1100 -1376 1165 -1359
rect 1378 -1376 1443 -1360
rect 1100 -1410 1115 -1376
rect 1149 -1410 1393 -1376
rect 1427 -1410 1443 -1376
rect 1100 -1426 1165 -1410
rect 1378 -1426 1443 -1410
rect 1115 -1448 1145 -1426
rect 1028 -1703 1058 -1648
<< polycont >>
rect 1115 -1410 1149 -1376
rect 1393 -1410 1427 -1376
<< locali >>
rect 982 -837 1172 -803
rect 982 -904 1016 -837
rect 1138 -931 1172 -837
rect 1138 -965 1303 -931
rect 982 -1333 1010 -1299
rect 1157 -1333 1303 -1299
rect 982 -1376 1016 -1333
rect 982 -1410 1115 -1376
rect 1149 -1410 1165 -1376
rect 982 -1444 1016 -1410
rect 982 -1478 1010 -1444
rect 1269 -1521 1303 -1333
rect 1377 -1410 1393 -1376
rect 1427 -1410 1443 -1376
rect 982 -1945 1016 -1903
rect 982 -1979 1270 -1945
<< viali >>
rect 1115 -1410 1149 -1376
rect 1393 -1410 1427 -1376
<< metal1 >>
rect 1315 -894 1381 -839
rect 1409 -950 1437 -935
rect 1064 -1056 1104 -1050
rect 1064 -1129 1110 -1056
rect 1269 -1193 1303 -1129
rect 1100 -1370 1165 -1369
rect 1100 -1376 1171 -1370
rect 1100 -1410 1115 -1376
rect 1149 -1410 1171 -1376
rect 1100 -1416 1171 -1410
rect 1268 -1448 1303 -1193
rect 1378 -1376 1449 -1369
rect 1378 -1410 1393 -1376
rect 1427 -1410 1449 -1376
rect 1378 -1416 1449 -1410
rect 1151 -1486 1303 -1448
rect 1151 -1494 1197 -1486
rect 1064 -1702 1110 -1648
rect 1419 -1975 1447 -1929
rect 1315 -2053 1391 -2007
use sky130_fd_pr__nfet_01v8_QRJQW7  M1
timestamp 1741451707
transform 1 0 1130 0 1 -1548
box -65 -126 73 126
use sky130_fd_pr__nfet_01v8_2SPF2Z  M2
timestamp 1741451707
transform 1 0 1043 0 1 -1802
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_2JZFD3  M3
timestamp 1741456812
transform 1 0 1043 0 1 -1517
box -73 -157 73 95
use sky130_fd_pr__pfet_01v8_EJJ636_2  M4
timestamp 1741452760
transform 1 0 1130 0 1 -1229
box -65 -136 153 162
use sky130_fd_pr__pfet_01v8_EJJ636  M5
timestamp 1741454074
transform 1 0 1043 0 1 -1229
box -109 -136 109 162
use sky130_fd_pr__pfet_01v8_WXG636  M6
timestamp 1741454074
transform 1 0 1043 0 1 -975
box -109 -136 109 136
use sky130_fd_pr__nfet_01v8_3RATTY  M88
timestamp 1741541561
transform 1 0 1355 0 1 -1781
box -98 -282 98 282
use sky130_fd_pr__pfet_01v8_HW9MHL  M99
timestamp 1741459568
transform 1 0 1350 0 1 -999
box -129 -198 129 160
<< end >>
