** sch_path: /foss/designs/tt10-uR-IPs/xschem/PTAT_wulff_tb.sch
**.subckt PTAT_wulff_tb
x1 in GND out PTAT_wulff
XR10 GND out GND sky130_fd_pr__res_xhigh_po_0p35 L=0.175 mult=1 m=1
E1 in GND VOL=' 1.8+(0.1*1.8*SIN(time*2*pi*1e6)) '
**** begin user architecture code


.param Vdd = 1.8V
.param V60Hz = 0.1

*V_PS_DC in GND {Vdd} DC
*V_PS_ripple in GND SIN(time*2*pi*1e6)

.control

*op
tran 10n 1u

write tb_ptat.raw

.endc



** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  PTAT_wulff.sym # of pins=3
** sym_path: /foss/designs/tt10-uR-IPs/xschem/PTAT_wulff.sym
** sch_path: /foss/designs/tt10-uR-IPs/xschem/PTAT_wulff.sch
.subckt PTAT_wulff Vdd Vss Iptat
*.ipin Vdd
*.ipin Vss
*.opin Iptat
XM10 Iptat Iptat Vdd Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 net1 net4 Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR10 net2 net3 Vss sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XD2 net1 Vss sky130_fd_pr__diode_pw2nd_11v0 area=1e12 perim=4e6
XD1 net2 Vss sky130_fd_pr__diode_pw2nd_11v0 area=1e12 perim=4e6
XM2 Vdd Iptat net4 Vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Iptat net1 net3 Vss sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
