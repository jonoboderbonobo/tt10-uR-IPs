magic
tech sky130A
magscale 1 2
timestamp 1738086101
<< checkpaint >>
rect 61 1605 3003 1658
rect 61 1552 3372 1605
rect 61 -1682 3741 1552
rect 430 -1735 3741 -1682
rect 799 -1788 3741 -1735
<< error_s >>
rect 485 1305 520 1339
rect 486 1286 520 1305
rect 294 1237 356 1243
rect 294 1203 306 1237
rect 294 1197 356 1203
rect 294 -91 356 -85
rect 294 -125 306 -91
rect 294 -131 356 -125
rect 505 -227 520 1286
rect 539 1252 574 1286
rect 894 1252 929 1286
rect 539 -227 573 1252
rect 895 1233 929 1252
rect 703 1184 765 1190
rect 703 1150 715 1184
rect 703 1144 765 1150
rect 703 -144 765 -138
rect 703 -178 715 -144
rect 703 -184 765 -178
rect 539 -261 554 -227
rect 914 -280 929 1233
rect 948 1199 983 1233
rect 948 -280 982 1199
rect 1112 1131 1174 1137
rect 1112 1097 1124 1131
rect 1112 1091 1174 1097
rect 1304 398 1338 416
rect 1304 362 1374 398
rect 1321 328 1392 362
rect 1672 328 1707 362
rect 1112 -197 1174 -191
rect 1112 -231 1124 -197
rect 1112 -237 1174 -231
rect 948 -314 963 -280
rect 1321 -333 1391 328
rect 1673 309 1707 328
rect 1503 260 1561 266
rect 1503 226 1515 260
rect 1503 220 1561 226
rect 1503 -250 1561 -244
rect 1503 -284 1515 -250
rect 1503 -290 1561 -284
rect 1321 -369 1374 -333
rect 1692 -386 1707 309
rect 1726 275 1761 309
rect 1726 -386 1760 275
rect 1872 207 1930 213
rect 1872 173 1884 207
rect 1872 167 1930 173
rect 1872 -303 1930 -297
rect 1872 -337 1884 -303
rect 1872 -343 1930 -337
rect 1726 -420 1741 -386
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM1
timestamp 0
transform 1 0 1901 0 1 -65
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM2
timestamp 0
transform 1 0 734 0 1 503
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM3
timestamp 0
transform 1 0 2270 0 1 -118
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM4
timestamp 0
transform 1 0 1143 0 1 450
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM6
timestamp 0
transform 1 0 1532 0 1 -12
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM10
timestamp 0
transform 1 0 325 0 1 556
box -231 -819 231 819
<< end >>
